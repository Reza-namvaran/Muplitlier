LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Multiplier_4x4 IS
    PORT (
        A : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        P : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
        -- Product term would have 8 bits;
    );
END Multiplier_4x4;

ARCHITECTURE BEHAVIORAL OF Multiplier_4x4 IS
BEGIN
    -- TODO
END BEHAVIORAL;
